library verilog;
use verilog.vl_types.all;
entity RALU_vlg_vec_tst is
end RALU_vlg_vec_tst;
