library verilog;
use verilog.vl_types.all;
entity MCD_vlg_vec_tst is
end MCD_vlg_vec_tst;
