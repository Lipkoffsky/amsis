library verilog;
use verilog.vl_types.all;
entity ALU_ParallelCarry_vlg_vec_tst is
end ALU_ParallelCarry_vlg_vec_tst;
